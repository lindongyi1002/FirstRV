/*==============================================================================================
    Filename            :   ALU.v
    Author              :   Lindongyi
    Description         :   1. 可以实现与或加减功能, 可以实现小于比较置位功能, 可以实现或非功能;
                            2. 使用4位输入控制ALU功能;
                            3. 纯组合逻辑电路; 
    Called by           :   
    Revision History    :   23-05-02
    Email               :   1292471097@qq.com
    Company             :   Jiang Group of Center for Carbon-based Electronics, Peking University
    Copyright           :   2023, Lindongyi, All right reserved
==============================================================================================*/

module ALU(

);
endmodule